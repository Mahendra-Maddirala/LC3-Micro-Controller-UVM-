//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: 
// This file contains defines and typedefs to be compiled for use in
// the simulation running on the emulator when using Veloce.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
                                                                               

typedef bit [1:0] mem_state_t;
typedef bit [15:0] DMem_addr_t;
typedef bit [15:0] DMem_din_t;
typedef bit DMem_rd_t;
typedef bit [15:0] memout_t;

// pragma uvmf custom additional begin
// pragma uvmf custom additional end

